library verilog;
use verilog.vl_types.all;
entity FinalTestBench is
end FinalTestBench;
