library verilog;
use verilog.vl_types.all;
entity invclass is
    port(
        a               : in     vl_logic;
        w               : out    vl_logic
    );
end invclass;
