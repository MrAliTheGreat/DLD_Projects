`timescale 1ns/1ns
module smbs_TB();
  reg serIn;
  reg [3:0] PB;
  reg [1:0] LB;
  reg [3:0][3:0] L;
  smbs cut_broadcaster (serIn, PB, LB, L);
  initial begin
    serIn = 1'b0;
    PB = 4'b0000;
    LB = 2'b00;
    #100;
    serIn = 1'b1;
    PB = 4'b0001;
    LB = 2'b10;
    #100;
    serIn = 1'b1;
    PB = 4'b0011;
    LB = 2'b01;
    #100;
    serIn = 1'b0;
    PB = 4'b1001;
    LB = 2'b11;
    #100;
    serIn = 1'b1;
    PB = 4'b0111;
    LB = 2'b01;
    #100;
    serIn = 1'b1;
    PB = 4'b1101;
    LB = 2'b10;
    #100;
    serIn = 1'b1;
    PB = 4'b1111;
    LB = 2'b11;
    #100;
    serIn = 1'b0;
    PB = 4'b0101;
    LB = 2'b10;
    #100;
    serIn = 1'b1;
    PB = 4'b1110;
    LB = 2'b00;
    #100;
    serIn = 1'b1;
    PB = 4'b0000;
    #100;
    serIn = 1'b1;
    PB = 4'b1100;
    #100;
    serIn = 1'b0;
    PB = 4'b1000;
    LB = 2'b10;
    #100;
    $stop;
  end
endmodule

module six_bit_shift_register_TB();
  logic clk;
  logic rst;
  logic en;
  logic serIn;
  logic [0:5]Q;
  six_bit_shift_register cut_Shift (serIn, clk, rst, en, Q);
  initial begin
    serIn = 1'b0;
    rst = 1'b0;
    en = 1'b1;
    clk = 1'b0;
    #100;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b0;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b0;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    $stop;
  end
endmodule

module sreg6_TB();
  logic clk;
  logic rst;
  logic en;
  logic serIn;
  logic [0:5]Q;
  SReg6 cut_sreg6 (clk, rst, en, serIn, Q);
  initial begin
    serIn = 1'b0;
    rst = 1'b0;
    en = 1'b1;
    clk = 1'b0;
    #100;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b0;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b1;
    clk = 1'b0;
    #100;
    serIn = 1'b1;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    serIn = 1'b0;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    clk = 1'b0;
    #100;
    serIn = 1'b0;
    clk = 1'b1;
    #100;
    $stop;
  end
endmodule
/*
module controller_TB();
logic in;
logic clk;
logic rst;
logic en;
logic port_en;
logic smbs_en;
logic out;
controller CUT (clk ,rst ,en, in ,out, port_en, smbs_en);
initial begin
  #100 in = 1;
  rst = 1'b0;
  en = 1'b1;
  #50 clk = 1;
  #50 clk = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 0;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50 in = 1;
  #50 clk = 1;
  #50 clk = 0;
  #50
  $stop;
  end
endmodule
*/
