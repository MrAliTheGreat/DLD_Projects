library verilog;
use verilog.vl_types.all;
entity sreg6_TB is
end sreg6_TB;
