library verilog;
use verilog.vl_types.all;
entity smbs_TB is
end smbs_TB;
