library verilog;
use verilog.vl_types.all;
entity demultiTB is
end demultiTB;
