library verilog;
use verilog.vl_types.all;
entity demultiplexer_4selectTB is
end demultiplexer_4selectTB;
