library verilog;
use verilog.vl_types.all;
entity Final_TestBench is
end Final_TestBench;
