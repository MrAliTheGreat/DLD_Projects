library verilog;
use verilog.vl_types.all;
entity input_wrapper_TB is
end input_wrapper_TB;
