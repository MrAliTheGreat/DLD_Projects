library verilog;
use verilog.vl_types.all;
entity controller_TB is
end controller_TB;
