library verilog;
use verilog.vl_types.all;
entity inv_nor2_3TB is
end inv_nor2_3TB;
