library verilog;
use verilog.vl_types.all;
entity demulti2TB is
end demulti2TB;
