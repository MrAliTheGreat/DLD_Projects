library verilog;
use verilog.vl_types.all;
entity demulti2_gateTB is
end demulti2_gateTB;
