library verilog;
use verilog.vl_types.all;
entity demulti4_gate_allTB is
end demulti4_gate_allTB;
