library verilog;
use verilog.vl_types.all;
entity DataPath_TB is
end DataPath_TB;
