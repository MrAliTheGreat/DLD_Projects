library verilog;
use verilog.vl_types.all;
entity demulti4TB is
end demulti4TB;
