library verilog;
use verilog.vl_types.all;
entity demultiplexer_2selectTB is
end demultiplexer_2selectTB;
