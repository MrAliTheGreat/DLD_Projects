library verilog;
use verilog.vl_types.all;
entity output_wrapper_TB is
end output_wrapper_TB;
