library verilog;
use verilog.vl_types.all;
entity demultiplexer4_selectTB is
end demultiplexer4_selectTB;
