library verilog;
use verilog.vl_types.all;
entity six_bit_shift_register_TB is
end six_bit_shift_register_TB;
