library verilog;
use verilog.vl_types.all;
entity broadcasterTB is
end broadcasterTB;
