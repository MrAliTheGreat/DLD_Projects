library verilog;
use verilog.vl_types.all;
entity demultiplexerTB is
end demultiplexerTB;
