module controller_TB();
  reg clk;
  reg rst;
  reg start;
  reg [7:0] y;
  reg signed [16:0] exp;
  
  wire ready , ldx , ldy , ldterm , ldexp , init_term , init_exp , minus1_en , x_en , i_en , iplus_en;
  wire [3:0] counteri , counteriplus;  
  Controller cut_controller(clk , rst , start , y , exp , ready , ldx , ldy , ldterm , ldexp , init_term , init_exp , minus1_en , x_en , i_en , iplus_en , counteri , counteriplus);
  initial begin
    #100;
    rst = 1;
    y = 8'b0_0001000;
    exp = 17'b000000000_00000010;
    start = 0;
    clk = 0;
    #50;
    rst = 0;
    start = 1;
    #10 clk = 1;
    #100 clk = 0;
    start = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #200
    $stop;
  end
endmodule


module DataPath_TB();
  reg clk;
  reg rst;
  reg start;
  reg signed [16:0] x;
  reg [7:0] y;
  
  wire ready;
  wire signed [16:0] Rout;
  Circuit cut_controller_and_circuit(clk , rst , start , x , y , ready , Rout);
  initial begin
    #100;
    rst = 1;
    y = 8'b0_0001000;
    x = 17'b000000000_00000010;
    start = 0;
    clk = 0;
    #50;
    rst = 0;
    start = 1;
    #10 clk = 1;
    #100 clk = 0;
    start = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #50 clk = 1;
    #50 clk = 0;
    #200
    $stop;
  end
endmodule


