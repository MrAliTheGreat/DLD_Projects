library verilog;
use verilog.vl_types.all;
entity line_seperator is
    port(
        L               : in     vl_logic_vector(3 downto 0);
        L0              : out    vl_logic;
        L1              : out    vl_logic;
        L2              : out    vl_logic;
        L3              : out    vl_logic;
        L4              : out    vl_logic;
        L5              : out    vl_logic;
        L6              : out    vl_logic;
        L7              : out    vl_logic;
        L8              : out    vl_logic;
        L9              : out    vl_logic;
        L10             : out    vl_logic;
        L11             : out    vl_logic;
        L12             : out    vl_logic;
        L13             : out    vl_logic;
        L14             : out    vl_logic;
        L15             : out    vl_logic
    );
end line_seperator;
