library verilog;
use verilog.vl_types.all;
entity demulti4_gateTB is
end demulti4_gateTB;
